library verilog;
use verilog.vl_types.all;
entity testbench4 is
end testbench4;

library verilog;
use verilog.vl_types.all;
entity testbench22 is
end testbench22;

library verilog;
use verilog.vl_types.all;
entity testbench2 is
end testbench2;

library verilog;
use verilog.vl_types.all;
entity testbench12 is
end testbench12;

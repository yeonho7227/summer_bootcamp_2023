library verilog;
use verilog.vl_types.all;
entity testbench3 is
end testbench3;

library verilog;
use verilog.vl_types.all;
entity testbench5 is
end testbench5;

library verilog;
use verilog.vl_types.all;
entity testbench9 is
end testbench9;

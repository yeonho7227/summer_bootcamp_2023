library verilog;
use verilog.vl_types.all;
entity testbench6 is
end testbench6;

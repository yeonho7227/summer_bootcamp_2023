library verilog;
use verilog.vl_types.all;
entity testbench11 is
end testbench11;
